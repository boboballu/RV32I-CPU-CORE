../fifo/fifo.sv