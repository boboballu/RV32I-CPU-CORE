// Author: Tarun Govind Kesavamurthi
// School: North Carolina State University
// mail  : tkesava@ncsu.edu
/********************************************************************************/
//debug_headerfile is instanced in all the files
// comment the definition below to disable debugging io at mem stage (mem_debug)
//`define mem_debug
//`define BR_RESOLVE_D
//`define BR_RESOLVE_M
/********************************************************************************/
// testbench.sv variables
int CONSOLE_ADDR = 65532;
int EXE_TIME	 = 20000;
/********************************************************************************/

