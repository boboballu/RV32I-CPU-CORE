// Author: Tarun Govind Kesavamurthi
// School: North Carolina State University
// mail  : tkesava@ncsu.edu
/********************************************************************************/
// comment the definition below to disable debugging io at mem stage (mem_debug)
`define mem_debug
//`define BR_RESOLVE_D
//`define BR_RESOLVE_M