../n_ff_cdc/sync.sv