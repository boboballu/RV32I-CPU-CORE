../skid_buffer/ready_valid_if.sv