
`define mem_debug

